// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// pcie_ed.v

// Generated using ACDS version 22.1 174

`timescale 1 ps / 1 ps
module pcie_ed (
		input  wire  hip_serial_rx_n_in0,   // hip_serial.rx_n_in0
		input  wire  hip_serial_rx_n_in1,   //           .rx_n_in1
		input  wire  hip_serial_rx_n_in2,   //           .rx_n_in2
		input  wire  hip_serial_rx_n_in3,   //           .rx_n_in3
		input  wire  hip_serial_rx_n_in4,   //           .rx_n_in4
		input  wire  hip_serial_rx_n_in5,   //           .rx_n_in5
		input  wire  hip_serial_rx_n_in6,   //           .rx_n_in6
		input  wire  hip_serial_rx_n_in7,   //           .rx_n_in7
		input  wire  hip_serial_rx_n_in8,   //           .rx_n_in8
		input  wire  hip_serial_rx_n_in9,   //           .rx_n_in9
		input  wire  hip_serial_rx_n_in10,  //           .rx_n_in10
		input  wire  hip_serial_rx_n_in11,  //           .rx_n_in11
		input  wire  hip_serial_rx_n_in12,  //           .rx_n_in12
		input  wire  hip_serial_rx_n_in13,  //           .rx_n_in13
		input  wire  hip_serial_rx_n_in14,  //           .rx_n_in14
		input  wire  hip_serial_rx_n_in15,  //           .rx_n_in15
		input  wire  hip_serial_rx_p_in0,   //           .rx_p_in0
		input  wire  hip_serial_rx_p_in1,   //           .rx_p_in1
		input  wire  hip_serial_rx_p_in2,   //           .rx_p_in2
		input  wire  hip_serial_rx_p_in3,   //           .rx_p_in3
		input  wire  hip_serial_rx_p_in4,   //           .rx_p_in4
		input  wire  hip_serial_rx_p_in5,   //           .rx_p_in5
		input  wire  hip_serial_rx_p_in6,   //           .rx_p_in6
		input  wire  hip_serial_rx_p_in7,   //           .rx_p_in7
		input  wire  hip_serial_rx_p_in8,   //           .rx_p_in8
		input  wire  hip_serial_rx_p_in9,   //           .rx_p_in9
		input  wire  hip_serial_rx_p_in10,  //           .rx_p_in10
		input  wire  hip_serial_rx_p_in11,  //           .rx_p_in11
		input  wire  hip_serial_rx_p_in12,  //           .rx_p_in12
		input  wire  hip_serial_rx_p_in13,  //           .rx_p_in13
		input  wire  hip_serial_rx_p_in14,  //           .rx_p_in14
		input  wire  hip_serial_rx_p_in15,  //           .rx_p_in15
		output wire  hip_serial_tx_n_out0,  //           .tx_n_out0
		output wire  hip_serial_tx_n_out1,  //           .tx_n_out1
		output wire  hip_serial_tx_n_out2,  //           .tx_n_out2
		output wire  hip_serial_tx_n_out3,  //           .tx_n_out3
		output wire  hip_serial_tx_n_out4,  //           .tx_n_out4
		output wire  hip_serial_tx_n_out5,  //           .tx_n_out5
		output wire  hip_serial_tx_n_out6,  //           .tx_n_out6
		output wire  hip_serial_tx_n_out7,  //           .tx_n_out7
		output wire  hip_serial_tx_n_out8,  //           .tx_n_out8
		output wire  hip_serial_tx_n_out9,  //           .tx_n_out9
		output wire  hip_serial_tx_n_out10, //           .tx_n_out10
		output wire  hip_serial_tx_n_out11, //           .tx_n_out11
		output wire  hip_serial_tx_n_out12, //           .tx_n_out12
		output wire  hip_serial_tx_n_out13, //           .tx_n_out13
		output wire  hip_serial_tx_n_out14, //           .tx_n_out14
		output wire  hip_serial_tx_n_out15, //           .tx_n_out15
		output wire  hip_serial_tx_p_out0,  //           .tx_p_out0
		output wire  hip_serial_tx_p_out1,  //           .tx_p_out1
		output wire  hip_serial_tx_p_out2,  //           .tx_p_out2
		output wire  hip_serial_tx_p_out3,  //           .tx_p_out3
		output wire  hip_serial_tx_p_out4,  //           .tx_p_out4
		output wire  hip_serial_tx_p_out5,  //           .tx_p_out5
		output wire  hip_serial_tx_p_out6,  //           .tx_p_out6
		output wire  hip_serial_tx_p_out7,  //           .tx_p_out7
		output wire  hip_serial_tx_p_out8,  //           .tx_p_out8
		output wire  hip_serial_tx_p_out9,  //           .tx_p_out9
		output wire  hip_serial_tx_p_out10, //           .tx_p_out10
		output wire  hip_serial_tx_p_out11, //           .tx_p_out11
		output wire  hip_serial_tx_p_out12, //           .tx_p_out12
		output wire  hip_serial_tx_p_out13, //           .tx_p_out13
		output wire  hip_serial_tx_p_out14, //           .tx_p_out14
		output wire  hip_serial_tx_p_out15, //           .tx_p_out15
		input  wire  refclk0_clk,           //    refclk0.clk
		input  wire  refclk1_clk,           //    refclk1.clk
		input  wire  pin_perst_reset_n      //  pin_perst.reset_n
	);

	wire           dut_p0_rx_st0_valid;                         // dut:p0_rx_st0_dvalid_o -> pio0:pio_rx_st0_dvalid_i
	wire   [255:0] dut_p0_rx_st0_data;                          // dut:p0_rx_st0_data_o -> pio0:pio_rx_st0_payload_i
	wire           dut_p0_rx_st0_ready;                         // pio0:pio_rx_st_ready_o -> dut:p0_rx_st_ready_i
	wire           dut_p0_rx_st0_startofpacket;                 // dut:p0_rx_st0_sop_o -> pio0:pio_rx_st0_sop_i
	wire           dut_p0_rx_st0_endofpacket;                   // dut:p0_rx_st0_eop_o -> pio0:pio_rx_st0_eop_i
	wire     [2:0] dut_p0_rx_st0_empty;                         // dut:p0_rx_st0_empty_o -> pio0:pio_rx_st0_empty_i
	wire           dut_p0_rx_st1_valid;                         // dut:p0_rx_st1_dvalid_o -> pio0:pio_rx_st1_dvalid_i
	wire   [255:0] dut_p0_rx_st1_data;                          // dut:p0_rx_st1_data_o -> pio0:pio_rx_st1_payload_i
	wire           dut_p0_rx_st1_startofpacket;                 // dut:p0_rx_st1_sop_o -> pio0:pio_rx_st1_sop_i
	wire           dut_p0_rx_st1_endofpacket;                   // dut:p0_rx_st1_eop_o -> pio0:pio_rx_st1_eop_i
	wire     [2:0] dut_p0_rx_st1_empty;                         // dut:p0_rx_st1_empty_o -> pio0:pio_rx_st1_empty_i
	wire           dut_p0_rx_st2_valid;                         // dut:p0_rx_st2_dvalid_o -> pio0:pio_rx_st2_dvalid_i
	wire   [255:0] dut_p0_rx_st2_data;                          // dut:p0_rx_st2_data_o -> pio0:pio_rx_st2_payload_i
	wire           dut_p0_rx_st2_startofpacket;                 // dut:p0_rx_st2_sop_o -> pio0:pio_rx_st2_sop_i
	wire           dut_p0_rx_st2_endofpacket;                   // dut:p0_rx_st2_eop_o -> pio0:pio_rx_st2_eop_i
	wire     [2:0] dut_p0_rx_st2_empty;                         // dut:p0_rx_st2_empty_o -> pio0:pio_rx_st2_empty_i
	wire           dut_p0_rx_st3_valid;                         // dut:p0_rx_st3_dvalid_o -> pio0:pio_rx_st3_dvalid_i
	wire   [255:0] dut_p0_rx_st3_data;                          // dut:p0_rx_st3_data_o -> pio0:pio_rx_st3_payload_i
	wire           dut_p0_rx_st3_startofpacket;                 // dut:p0_rx_st3_sop_o -> pio0:pio_rx_st3_sop_i
	wire           dut_p0_rx_st3_endofpacket;                   // dut:p0_rx_st3_eop_o -> pio0:pio_rx_st3_eop_i
	wire     [2:0] dut_p0_rx_st3_empty;                         // dut:p0_rx_st3_empty_o -> pio0:pio_rx_st3_empty_i
	wire           pio0_tx_st0_pio_valid;                       // pio0:pio_tx_st0_dvalid_o -> dut:p0_tx_st0_dvalid_i
	wire   [255:0] pio0_tx_st0_pio_data;                        // pio0:pio_tx_st0_payload_o -> dut:p0_tx_st0_data_i
	wire           pio0_tx_st0_pio_ready;                       // dut:p0_tx_st_ready_o -> pio0:pio_tx_st_ready_i
	wire           pio0_tx_st0_pio_startofpacket;               // pio0:pio_tx_st0_sop_o -> dut:p0_tx_st0_sop_i
	wire           pio0_tx_st0_pio_endofpacket;                 // pio0:pio_tx_st0_eop_o -> dut:p0_tx_st0_eop_i
	wire           pio0_tx_st1_pio_valid;                       // pio0:pio_tx_st1_dvalid_o -> dut:p0_tx_st1_dvalid_i
	wire   [255:0] pio0_tx_st1_pio_data;                        // pio0:pio_tx_st1_payload_o -> dut:p0_tx_st1_data_i
	wire           pio0_tx_st1_pio_startofpacket;               // pio0:pio_tx_st1_sop_o -> dut:p0_tx_st1_sop_i
	wire           pio0_tx_st1_pio_endofpacket;                 // pio0:pio_tx_st1_eop_o -> dut:p0_tx_st1_eop_i
	wire           pio0_tx_st2_pio_valid;                       // pio0:pio_tx_st2_dvalid_o -> dut:p0_tx_st2_dvalid_i
	wire   [255:0] pio0_tx_st2_pio_data;                        // pio0:pio_tx_st2_payload_o -> dut:p0_tx_st2_data_i
	wire           pio0_tx_st2_pio_startofpacket;               // pio0:pio_tx_st2_sop_o -> dut:p0_tx_st2_sop_i
	wire           pio0_tx_st2_pio_endofpacket;                 // pio0:pio_tx_st2_eop_o -> dut:p0_tx_st2_eop_i
	wire           pio0_tx_st3_pio_valid;                       // pio0:pio_tx_st3_dvalid_o -> dut:p0_tx_st3_dvalid_i
	wire   [255:0] pio0_tx_st3_pio_data;                        // pio0:pio_tx_st3_payload_o -> dut:p0_tx_st3_data_i
	wire           pio0_tx_st3_pio_startofpacket;               // pio0:pio_tx_st3_sop_o -> dut:p0_tx_st3_sop_i
	wire           pio0_tx_st3_pio_endofpacket;                 // pio0:pio_tx_st3_eop_o -> dut:p0_tx_st3_eop_i
	wire           dut_coreclkout_hip_clk;                      // dut:coreclkout_hip -> pio0:Clk_i
	wire           pio0_pio_master_clk_clk;                     // pio0:pio_clk -> [MEM0:clk, mm_interconnect_0:pio0_pio_master_clk_clk, rst_controller:clk]
	wire    [31:0] dut_p0_rx_st_misc_rx_st1_prefix;             // dut:p0_rx_st1_prefix_o -> pio0:pio_rx_st1_tlp_prfx_i
	wire           dut_p0_rx_st_misc_rx_st2_pvalid;             // dut:p0_rx_st2_pvalid_o -> pio0:pio_rx_st2_pvalid_i
	wire    [31:0] dut_p0_rx_st_misc_rx_st0_prefix;             // dut:p0_rx_st0_prefix_o -> pio0:pio_rx_st0_tlp_prfx_i
	wire   [127:0] dut_p0_rx_st_misc_rx_st3_hdr;                // dut:p0_rx_st3_hdr_o -> pio0:pio_rx_st3_header_i
	wire           dut_p0_rx_st_misc_rx_st0_pvalid;             // dut:p0_rx_st0_pvalid_o -> pio0:pio_rx_st0_pvalid_i
	wire           dut_p0_rx_st_misc_rx_st1_pvalid;             // dut:p0_rx_st1_pvalid_o -> pio0:pio_rx_st1_pvalid_i
	wire    [31:0] dut_p0_rx_st_misc_rx_st2_prefix;             // dut:p0_rx_st2_prefix_o -> pio0:pio_rx_st2_tlp_prfx_i
	wire    [31:0] dut_p0_rx_st_misc_rx_st3_prefix;             // dut:p0_rx_st3_prefix_o -> pio0:pio_rx_st3_tlp_prfx_i
	wire           dut_p0_rx_st_misc_rx_st3_pvalid;             // dut:p0_rx_st3_pvalid_o -> pio0:pio_rx_st3_pvalid_i
	wire   [127:0] dut_p0_rx_st_misc_rx_st2_hdr;                // dut:p0_rx_st2_hdr_o -> pio0:pio_rx_st2_header_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st0_bar;                // dut:p0_rx_st0_bar_o -> pio0:pio_rx_st0_bar_i
	wire     [2:0] pio0_rx_st0_pio_misc_rx_st_dcrdt_init;       // pio0:rx_st_dcrdt_init_o -> dut:p0_rx_st_dcrdt_init_i
	wire     [2:0] pio0_rx_st0_pio_misc_rx_st_hcrdt_update;     // pio0:rx_st_hcrdt_update_o -> dut:p0_rx_st_hcrdt_update_i
	wire    [11:0] pio0_rx_st0_pio_misc_rx_st_dcrdt_update_cnt; // pio0:rx_st_dcrdt_update_cnt_o -> dut:p0_rx_st_dcrdt_update_cnt_i
	wire     [2:0] pio0_rx_st0_pio_misc_rx_st_dcrdt_update;     // pio0:rx_st_dcrdt_update_o -> dut:p0_rx_st_dcrdt_update_i
	wire     [5:0] pio0_rx_st0_pio_misc_rx_st_hcrdt_update_cnt; // pio0:rx_st_hcrdt_update_cnt_o -> dut:p0_rx_st_hcrdt_update_cnt_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st1_bar;                // dut:p0_rx_st1_bar_o -> pio0:pio_rx_st1_bar_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st_hcrdt_init_ack;      // dut:p0_rx_st_hcrdt_init_ack_o -> pio0:rx_st_hcrdt_init_ack_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st_dcrdt_init_ack;      // dut:p0_rx_st_dcrdt_init_ack_o -> pio0:rx_st_dcrdt_init_ack_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st2_bar;                // dut:p0_rx_st2_bar_o -> pio0:pio_rx_st2_bar_i
	wire     [2:0] pio0_rx_st0_pio_misc_rx_st_hcrdt_init;       // pio0:rx_st_hcrdt_init_o -> dut:p0_rx_st_hcrdt_init_i
	wire   [127:0] dut_p0_rx_st_misc_rx_st0_hdr;                // dut:p0_rx_st0_hdr_o -> pio0:pio_rx_st0_header_i
	wire           dut_p0_rx_st_misc_rx_st0_hvalid;             // dut:p0_rx_st0_hvalid_o -> pio0:pio_rx_st0_hvalid_i
	wire           dut_p0_rx_st_misc_rx_st1_hvalid;             // dut:p0_rx_st1_hvalid_o -> pio0:pio_rx_st1_hvalid_i
	wire           dut_p0_rx_st_misc_rx_st2_hvalid;             // dut:p0_rx_st2_hvalid_o -> pio0:pio_rx_st2_hvalid_i
	wire           dut_p0_rx_st_misc_rx_st3_hvalid;             // dut:p0_rx_st3_hvalid_o -> pio0:pio_rx_st3_hvalid_i
	wire   [127:0] dut_p0_rx_st_misc_rx_st1_hdr;                // dut:p0_rx_st1_hdr_o -> pio0:pio_rx_st1_header_i
	wire     [2:0] dut_p0_rx_st_misc_rx_st3_bar;                // dut:p0_rx_st3_bar_o -> pio0:pio_rx_st3_bar_i
	wire     [2:0] dut_p0_tx_st_misc_tx_st_hcrdt_init;          // dut:p0_tx_st_hcrdt_init_o -> pio0:tx_st_hcrdt_init_i
	wire           pio0_tx_st0_pio_misc_tx_st0_pvalid;          // pio0:pio_tx_st0_pvalid_o -> dut:p0_tx_st0_pvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st1_pvalid;          // pio0:pio_tx_st1_pvalid_o -> dut:p0_tx_st1_pvalid_i
	wire    [11:0] dut_p0_tx_st_misc_tx_st_dcrdt_update_cnt;    // dut:p0_tx_st_dcrdt_update_cnt_o -> pio0:tx_st_dcrdt_update_cnt_i
	wire   [127:0] pio0_tx_st0_pio_misc_tx_st1_hdr;             // pio0:pio_tx_st1_header_o -> dut:p0_tx_st1_hdr_i
	wire     [2:0] dut_p0_tx_st_misc_tx_st_dcrdt_init;          // dut:p0_tx_st_dcrdt_init_o -> pio0:tx_st_dcrdt_init_i
	wire   [127:0] pio0_tx_st0_pio_misc_tx_st3_hdr;             // pio0:pio_tx_st3_header_o -> dut:p0_tx_st3_hdr_i
	wire           pio0_tx_st0_pio_misc_tx_st2_pvalid;          // pio0:pio_tx_st2_pvalid_o -> dut:p0_tx_st2_pvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st3_pvalid;          // pio0:pio_tx_st3_pvalid_o -> dut:p0_tx_st3_pvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st1_hvalid;          // pio0:pio_tx_st1_hvalid_o -> dut:p0_tx_st1_hvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st2_hvalid;          // pio0:pio_tx_st2_hvalid_o -> dut:p0_tx_st2_hvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st3_hvalid;          // pio0:pio_tx_st3_hvalid_o -> dut:p0_tx_st3_hvalid_i
	wire           pio0_tx_st0_pio_misc_tx_st0_hvalid;          // pio0:pio_tx_st0_hvalid_o -> dut:p0_tx_st0_hvalid_i
	wire   [127:0] pio0_tx_st0_pio_misc_tx_st0_hdr;             // pio0:pio_tx_st0_header_o -> dut:p0_tx_st0_hdr_i
	wire     [5:0] dut_p0_tx_st_misc_tx_st_hcrdt_update_cnt;    // dut:p0_tx_st_hcrdt_update_cnt_o -> pio0:tx_st_hcrdt_update_cnt_i
	wire     [2:0] pio0_tx_st0_pio_misc_tx_st_dcrdt_init_ack;   // pio0:tx_st_dcrdt_init_ack_o -> dut:p0_tx_st_dcrdt_init_ack_i
	wire    [31:0] pio0_tx_st0_pio_misc_tx_st2_prefix;          // pio0:pio_tx_st2_prefix_o -> dut:p0_tx_st2_prefix_i
	wire    [31:0] pio0_tx_st0_pio_misc_tx_st3_prefix;          // pio0:pio_tx_st3_prefix_o -> dut:p0_tx_st3_prefix_i
	wire   [127:0] pio0_tx_st0_pio_misc_tx_st2_hdr;             // pio0:pio_tx_st2_header_o -> dut:p0_tx_st2_hdr_i
	wire     [2:0] pio0_tx_st0_pio_misc_tx_st_hcrdtt_init_ack;  // pio0:tx_st_hcrdt_init_ack_o -> dut:p0_tx_st_hcrdt_init_ack_i
	wire     [2:0] dut_p0_tx_st_misc_tx_st_dcrdt_update;        // dut:p0_tx_st_dcrdt_update_o -> pio0:tx_st_dcrdt_update_i
	wire    [31:0] pio0_tx_st0_pio_misc_tx_st0_prefix;          // pio0:pio_tx_st0_prefix_o -> dut:p0_tx_st0_prefix_i
	wire    [31:0] pio0_tx_st0_pio_misc_tx_st1_prefix;          // pio0:pio_tx_st1_prefix_o -> dut:p0_tx_st1_prefix_i
	wire     [2:0] dut_p0_tx_st_misc_tx_st_hcrdt_update;        // dut:p0_tx_st_hcrdt_update_o -> pio0:tx_st_hcrdt_update_i
	wire           resetip_ninit_done_reset;                    // resetIP:ninit_done -> dut:ninit_done
	wire           dut_p0_reset_status_n_reset;                 // dut:p0_reset_status_n -> pio0:Rstn_i
	wire           pio0_pio_master_reset_reset;                 // pio0:pio_rst_n -> [MEM0:reset, rst_controller:reset_in0]
	wire  [1023:0] pio0_pio_master_readdata;                    // mm_interconnect_0:pio0_pio_master_readdata -> pio0:pio_readdata_i
	wire           pio0_pio_master_waitrequest;                 // mm_interconnect_0:pio0_pio_master_waitrequest -> pio0:pio_waitrequest_i
	wire    [63:0] pio0_pio_master_address;                     // pio0:pio_address_o -> mm_interconnect_0:pio0_pio_master_address
	wire           pio0_pio_master_read;                        // pio0:pio_read_o -> mm_interconnect_0:pio0_pio_master_read
	wire   [127:0] pio0_pio_master_byteenable;                  // pio0:pio_byteenable_o -> mm_interconnect_0:pio0_pio_master_byteenable
	wire           pio0_pio_master_readdatavalid;               // mm_interconnect_0:pio0_pio_master_readdatavalid -> pio0:pio_readdatavalid_i
	wire     [1:0] pio0_pio_master_response;                    // mm_interconnect_0:pio0_pio_master_response -> pio0:pio_response_i
	wire           pio0_pio_master_write;                       // pio0:pio_write_o -> mm_interconnect_0:pio0_pio_master_write
	wire  [1023:0] pio0_pio_master_writedata;                   // pio0:pio_writedata_o -> mm_interconnect_0:pio0_pio_master_writedata
	wire     [3:0] pio0_pio_master_burstcount;                  // pio0:pio_burstcount_o -> mm_interconnect_0:pio0_pio_master_burstcount
	wire           mm_interconnect_0_mem0_s1_chipselect;        // mm_interconnect_0:MEM0_s1_chipselect -> MEM0:chipselect
	wire  [1023:0] mm_interconnect_0_mem0_s1_readdata;          // MEM0:readdata -> mm_interconnect_0:MEM0_s1_readdata
	wire     [7:0] mm_interconnect_0_mem0_s1_address;           // mm_interconnect_0:MEM0_s1_address -> MEM0:address
	wire   [127:0] mm_interconnect_0_mem0_s1_byteenable;        // mm_interconnect_0:MEM0_s1_byteenable -> MEM0:byteenable
	wire           mm_interconnect_0_mem0_s1_write;             // mm_interconnect_0:MEM0_s1_write -> MEM0:write
	wire  [1023:0] mm_interconnect_0_mem0_s1_writedata;         // mm_interconnect_0:MEM0_s1_writedata -> MEM0:writedata
	wire           mm_interconnect_0_mem0_s1_clken;             // mm_interconnect_0:MEM0_s1_clken -> MEM0:clken
	wire           rst_controller_reset_out_reset;              // rst_controller:reset_out -> [mm_interconnect_0:MEM0_reset1_reset_bridge_in_reset_reset, mm_interconnect_0:pio0_pio_master_translator_reset_reset_bridge_in_reset_reset]

	pcie_ed_MEM0 mem0 (
		.clk        (pio0_pio_master_clk_clk),              //   input,     width = 1,   clk1.clk
		.address    (mm_interconnect_0_mem0_s1_address),    //   input,     width = 8,     s1.address
		.clken      (mm_interconnect_0_mem0_s1_clken),      //   input,     width = 1,       .clken
		.chipselect (mm_interconnect_0_mem0_s1_chipselect), //   input,     width = 1,       .chipselect
		.write      (mm_interconnect_0_mem0_s1_write),      //   input,     width = 1,       .write
		.readdata   (mm_interconnect_0_mem0_s1_readdata),   //  output,  width = 1024,       .readdata
		.writedata  (mm_interconnect_0_mem0_s1_writedata),  //   input,  width = 1024,       .writedata
		.byteenable (mm_interconnect_0_mem0_s1_byteenable), //   input,   width = 128,       .byteenable
		.reset      (~pio0_pio_master_reset_reset)          //   input,     width = 1, reset1.reset
	);

/*	pcie_ed_dut dut (
		.p0_rx_st_ready_i             (dut_p0_rx_st0_ready),                         //   input,    width = 1,              p0_rx_st0.ready
		.p0_rx_st0_data_o             (dut_p0_rx_st0_data),                          //  output,  width = 256,                       .data
		.p0_rx_st0_sop_o              (dut_p0_rx_st0_startofpacket),                 //  output,    width = 1,                       .startofpacket
		.p0_rx_st0_eop_o              (dut_p0_rx_st0_endofpacket),                   //  output,    width = 1,                       .endofpacket
		.p0_rx_st0_dvalid_o           (dut_p0_rx_st0_valid),                         //  output,    width = 1,                       .valid
		.p0_rx_st0_empty_o            (dut_p0_rx_st0_empty),                         //  output,    width = 3,                       .empty
		.p0_rx_st0_hdr_o              (dut_p0_rx_st_misc_rx_st0_hdr),                //  output,  width = 128,          p0_rx_st_misc.rx_st0_hdr
		.p0_rx_st0_prefix_o           (dut_p0_rx_st_misc_rx_st0_prefix),             //  output,   width = 32,                       .rx_st0_prefix
		.p0_rx_st0_hvalid_o           (dut_p0_rx_st_misc_rx_st0_hvalid),             //  output,    width = 1,                       .rx_st0_hvalid
		.p0_rx_st0_pvalid_o           (dut_p0_rx_st_misc_rx_st0_pvalid),             //  output,    width = 1,                       .rx_st0_pvalid
		.p0_rx_st0_bar_o              (dut_p0_rx_st_misc_rx_st0_bar),                //  output,    width = 3,                       .rx_st0_bar
		.p0_rx_st0_pt_parity_o        (),                                            //  output,    width = 1,                       .rx_st0_pt_parity
		.p0_rx_st1_hdr_o              (dut_p0_rx_st_misc_rx_st1_hdr),                //  output,  width = 128,                       .rx_st1_hdr
		.p0_rx_st1_prefix_o           (dut_p0_rx_st_misc_rx_st1_prefix),             //  output,   width = 32,                       .rx_st1_prefix
		.p0_rx_st1_hvalid_o           (dut_p0_rx_st_misc_rx_st1_hvalid),             //  output,    width = 1,                       .rx_st1_hvalid
		.p0_rx_st1_pvalid_o           (dut_p0_rx_st_misc_rx_st1_pvalid),             //  output,    width = 1,                       .rx_st1_pvalid
		.p0_rx_st1_bar_o              (dut_p0_rx_st_misc_rx_st1_bar),                //  output,    width = 3,                       .rx_st1_bar
		.p0_rx_st1_pt_parity_o        (),                                            //  output,    width = 1,                       .rx_st1_pt_parity
		.p0_rx_st2_hdr_o              (dut_p0_rx_st_misc_rx_st2_hdr),                //  output,  width = 128,                       .rx_st2_hdr
		.p0_rx_st2_prefix_o           (dut_p0_rx_st_misc_rx_st2_prefix),             //  output,   width = 32,                       .rx_st2_prefix
		.p0_rx_st2_hvalid_o           (dut_p0_rx_st_misc_rx_st2_hvalid),             //  output,    width = 1,                       .rx_st2_hvalid
		.p0_rx_st2_pvalid_o           (dut_p0_rx_st_misc_rx_st2_pvalid),             //  output,    width = 1,                       .rx_st2_pvalid
		.p0_rx_st2_bar_o              (dut_p0_rx_st_misc_rx_st2_bar),                //  output,    width = 3,                       .rx_st2_bar
		.p0_rx_st2_pt_parity_o        (),                                            //  output,    width = 1,                       .rx_st2_pt_parity
		.p0_rx_st3_hdr_o              (dut_p0_rx_st_misc_rx_st3_hdr),                //  output,  width = 128,                       .rx_st3_hdr
		.p0_rx_st3_prefix_o           (dut_p0_rx_st_misc_rx_st3_prefix),             //  output,   width = 32,                       .rx_st3_prefix
		.p0_rx_st3_hvalid_o           (dut_p0_rx_st_misc_rx_st3_hvalid),             //  output,    width = 1,                       .rx_st3_hvalid
		.p0_rx_st3_pvalid_o           (dut_p0_rx_st_misc_rx_st3_pvalid),             //  output,    width = 1,                       .rx_st3_pvalid
		.p0_rx_st3_bar_o              (dut_p0_rx_st_misc_rx_st3_bar),                //  output,    width = 3,                       .rx_st3_bar
		.p0_rx_st3_pt_parity_o        (),                                            //  output,    width = 1,                       .rx_st3_pt_parity
		.p0_rx_st_hcrdt_init_i        (pio0_rx_st0_pio_misc_rx_st_hcrdt_init),       //   input,    width = 3,                       .rx_st_Hcrdt_init
		.p0_rx_st_hcrdt_update_i      (pio0_rx_st0_pio_misc_rx_st_hcrdt_update),     //   input,    width = 3,                       .rx_st_Hcrdt_update
		.p0_rx_st_hcrdt_update_cnt_i  (pio0_rx_st0_pio_misc_rx_st_hcrdt_update_cnt), //   input,    width = 6,                       .rx_st_Hcrdt_update_cnt
		.p0_rx_st_hcrdt_init_ack_o    (dut_p0_rx_st_misc_rx_st_hcrdt_init_ack),      //  output,    width = 3,                       .rx_st_Hcrdt_init_ack
		.p0_rx_st_dcrdt_init_i        (pio0_rx_st0_pio_misc_rx_st_dcrdt_init),       //   input,    width = 3,                       .rx_st_Dcrdt_init
		.p0_rx_st_dcrdt_update_i      (pio0_rx_st0_pio_misc_rx_st_dcrdt_update),     //   input,    width = 3,                       .rx_st_Dcrdt_update
		.p0_rx_st_dcrdt_update_cnt_i  (pio0_rx_st0_pio_misc_rx_st_dcrdt_update_cnt), //   input,   width = 12,                       .rx_st_Dcrdt_update_cnt
		.p0_rx_st_dcrdt_init_ack_o    (dut_p0_rx_st_misc_rx_st_dcrdt_init_ack),      //  output,    width = 3,                       .rx_st_Dcrdt_init_ack
		.p0_rx_st1_data_o             (dut_p0_rx_st1_data),                          //  output,  width = 256,              p0_rx_st1.data
		.p0_rx_st1_sop_o              (dut_p0_rx_st1_startofpacket),                 //  output,    width = 1,                       .startofpacket
		.p0_rx_st1_eop_o              (dut_p0_rx_st1_endofpacket),                   //  output,    width = 1,                       .endofpacket
		.p0_rx_st1_dvalid_o           (dut_p0_rx_st1_valid),                         //  output,    width = 1,                       .valid
		.p0_rx_st1_empty_o            (dut_p0_rx_st1_empty),                         //  output,    width = 3,                       .empty
		.p0_rx_st2_data_o             (dut_p0_rx_st2_data),                          //  output,  width = 256,              p0_rx_st2.data
		.p0_rx_st2_sop_o              (dut_p0_rx_st2_startofpacket),                 //  output,    width = 1,                       .startofpacket
		.p0_rx_st2_eop_o              (dut_p0_rx_st2_endofpacket),                   //  output,    width = 1,                       .endofpacket
		.p0_rx_st2_dvalid_o           (dut_p0_rx_st2_valid),                         //  output,    width = 1,                       .valid
		.p0_rx_st2_empty_o            (dut_p0_rx_st2_empty),                         //  output,    width = 3,                       .empty
		.p0_rx_st3_data_o             (dut_p0_rx_st3_data),                          //  output,  width = 256,              p0_rx_st3.data
		.p0_rx_st3_sop_o              (dut_p0_rx_st3_startofpacket),                 //  output,    width = 1,                       .startofpacket
		.p0_rx_st3_eop_o              (dut_p0_rx_st3_endofpacket),                   //  output,    width = 1,                       .endofpacket
		.p0_rx_st3_dvalid_o           (dut_p0_rx_st3_valid),                         //  output,    width = 1,                       .valid
		.p0_rx_st3_empty_o            (dut_p0_rx_st3_empty),                         //  output,    width = 3,                       .empty
		.p0_tx_st_hcrdt_init_o        (dut_p0_tx_st_misc_tx_st_hcrdt_init),          //  output,    width = 3,          p0_tx_st_misc.tx_st_Hcrdt_init
		.p0_tx_st_hcrdt_update_o      (dut_p0_tx_st_misc_tx_st_hcrdt_update),        //  output,    width = 3,                       .tx_st_Hcrdt_update
		.p0_tx_st_hcrdt_update_cnt_o  (dut_p0_tx_st_misc_tx_st_hcrdt_update_cnt),    //  output,    width = 6,                       .tx_st_Hcrdt_update_cnt
		.p0_tx_st_hcrdt_init_ack_i    (pio0_tx_st0_pio_misc_tx_st_hcrdtt_init_ack),  //   input,    width = 3,                       .tx_st_Hcrdtt_init_ack
		.p0_tx_st_dcrdt_init_o        (dut_p0_tx_st_misc_tx_st_dcrdt_init),          //  output,    width = 3,                       .tx_st_Dcrdt_init
		.p0_tx_st_dcrdt_update_o      (dut_p0_tx_st_misc_tx_st_dcrdt_update),        //  output,    width = 3,                       .tx_st_Dcrdt_update
		.p0_tx_st_dcrdt_update_cnt_o  (dut_p0_tx_st_misc_tx_st_dcrdt_update_cnt),    //  output,   width = 12,                       .tx_st_Dcrdt_update_cnt
		.p0_tx_st_dcrdt_init_ack_i    (pio0_tx_st0_pio_misc_tx_st_dcrdt_init_ack),   //   input,    width = 3,                       .tx_st_Dcrdt_init_ack
		.p0_tx_st0_hdr_i              (pio0_tx_st0_pio_misc_tx_st0_hdr),             //   input,  width = 128,                       .tx_st0_hdr
		.p0_tx_st0_prefix_i           (pio0_tx_st0_pio_misc_tx_st0_prefix),          //   input,   width = 32,                       .tx_st0_prefix
		.p0_tx_st0_hvalid_i           (pio0_tx_st0_pio_misc_tx_st0_hvalid),          //   input,    width = 1,                       .tx_st0_hvalid
		.p0_tx_st0_pvalid_i           (pio0_tx_st0_pio_misc_tx_st0_pvalid),          //   input,    width = 1,                       .tx_st0_pvalid
		.p0_tx_st1_hdr_i              (pio0_tx_st0_pio_misc_tx_st1_hdr),             //   input,  width = 128,                       .tx_st1_hdr
		.p0_tx_st1_prefix_i           (pio0_tx_st0_pio_misc_tx_st1_prefix),          //   input,   width = 32,                       .tx_st1_prefix
		.p0_tx_st1_hvalid_i           (pio0_tx_st0_pio_misc_tx_st1_hvalid),          //   input,    width = 1,                       .tx_st1_hvalid
		.p0_tx_st1_pvalid_i           (pio0_tx_st0_pio_misc_tx_st1_pvalid),          //   input,    width = 1,                       .tx_st1_pvalid
		.p0_tx_st2_hdr_i              (pio0_tx_st0_pio_misc_tx_st2_hdr),             //   input,  width = 128,                       .tx_st2_hdr
		.p0_tx_st2_prefix_i           (pio0_tx_st0_pio_misc_tx_st2_prefix),          //   input,   width = 32,                       .tx_st2_prefix
		.p0_tx_st2_hvalid_i           (pio0_tx_st0_pio_misc_tx_st2_hvalid),          //   input,    width = 1,                       .tx_st2_hvalid
		.p0_tx_st2_pvalid_i           (pio0_tx_st0_pio_misc_tx_st2_pvalid),          //   input,    width = 1,                       .tx_st2_pvalid
		.p0_tx_st3_hdr_i              (pio0_tx_st0_pio_misc_tx_st3_hdr),             //   input,  width = 128,                       .tx_st3_hdr
		.p0_tx_st3_prefix_i           (pio0_tx_st0_pio_misc_tx_st3_prefix),          //   input,   width = 32,                       .tx_st3_prefix
		.p0_tx_st3_hvalid_i           (pio0_tx_st0_pio_misc_tx_st3_hvalid),          //   input,    width = 1,                       .tx_st3_hvalid
		.p0_tx_st3_pvalid_i           (pio0_tx_st0_pio_misc_tx_st3_pvalid),          //   input,    width = 1,                       .tx_st3_pvalid
		.p0_tx_st_ready_o             (pio0_tx_st0_pio_ready),                       //  output,    width = 1,              p0_tx_st0.ready
		.p0_tx_st0_data_i             (pio0_tx_st0_pio_data),                        //   input,  width = 256,                       .data
		.p0_tx_st0_sop_i              (pio0_tx_st0_pio_startofpacket),               //   input,    width = 1,                       .startofpacket
		.p0_tx_st0_eop_i              (pio0_tx_st0_pio_endofpacket),                 //   input,    width = 1,                       .endofpacket
		.p0_tx_st0_dvalid_i           (pio0_tx_st0_pio_valid),                       //   input,    width = 1,                       .valid
		.p0_tx_st1_data_i             (pio0_tx_st1_pio_data),                        //   input,  width = 256,              p0_tx_st1.data
		.p0_tx_st1_sop_i              (pio0_tx_st1_pio_startofpacket),               //   input,    width = 1,                       .startofpacket
		.p0_tx_st1_eop_i              (pio0_tx_st1_pio_endofpacket),                 //   input,    width = 1,                       .endofpacket
		.p0_tx_st1_dvalid_i           (pio0_tx_st1_pio_valid),                       //   input,    width = 1,                       .valid
		.p0_tx_st2_data_i             (pio0_tx_st2_pio_data),                        //   input,  width = 256,              p0_tx_st2.data
		.p0_tx_st2_sop_i              (pio0_tx_st2_pio_startofpacket),               //   input,    width = 1,                       .startofpacket
		.p0_tx_st2_eop_i              (pio0_tx_st2_pio_endofpacket),                 //   input,    width = 1,                       .endofpacket
		.p0_tx_st2_dvalid_i           (pio0_tx_st2_pio_valid),                       //   input,    width = 1,                       .valid
		.p0_tx_st3_data_i             (pio0_tx_st3_pio_data),                        //   input,  width = 256,              p0_tx_st3.data
		.p0_tx_st3_sop_i              (pio0_tx_st3_pio_startofpacket),               //   input,    width = 1,                       .startofpacket
		.p0_tx_st3_eop_i              (pio0_tx_st3_pio_endofpacket),                 //   input,    width = 1,                       .endofpacket
		.p0_tx_st3_dvalid_i           (pio0_tx_st3_pio_valid),                       //   input,    width = 1,                       .valid
		.p0_tx_ehp_deallocate_empty_o (),                                            //  output,    width = 1,              p0_tx_ehp.tx_ehp_deallocate_empty
		.p0_reset_status_n            (dut_p0_reset_status_n_reset),                 //  output,    width = 1,      p0_reset_status_n.reset_n
		.p0_slow_reset_status_n       (),                                            //  output,    width = 1, p0_slow_reset_status_n.reset_n
		.p0_link_up_o                 (),                                            //  output,    width = 1,          p0_hip_status.link_up
		.p0_dl_up_o                   (),                                            //  output,    width = 1,                       .dl_up
		.p0_surprise_down_err_o       (),                                            //  output,    width = 1,                       .surprise_down_err
		.p0_dl_timer_update_o         (),                                            //  output,    width = 1,                       .dl_timer_update
		.p0_ltssm_state_delay_o       (),                                            //  output,    width = 6,                       .ltssm_state_delay
		.p0_ltssm_st_hipfifo_ovrflw_o (),                                            //  output,    width = 1,                       .ltssm_st_hipfifo_ovrflw
		.p0_app_xfer_pending_i        (),                                            //   input,    width = 1,          p0_power_mgnt.app_xfer_pending
		.p0_pld_gp_status_i           (),                                            //   input,    width = 8,              p0_pld_gp.status
		.p0_pld_gp_ctrl_o             (),                                            //  output,    width = 8,                       .ctrl
		.p0_pld_gp_status_ready_o     (),                                            //  output,    width = 1,                       .status_ready
		.rx_n_in0                     (hip_serial_rx_n_in0),                         //   input,    width = 1,             hip_serial.rx_n_in0
		.rx_n_in1                     (hip_serial_rx_n_in1),                         //   input,    width = 1,                       .rx_n_in1
		.rx_n_in2                     (hip_serial_rx_n_in2),                         //   input,    width = 1,                       .rx_n_in2
		.rx_n_in3                     (hip_serial_rx_n_in3),                         //   input,    width = 1,                       .rx_n_in3
		.rx_n_in4                     (hip_serial_rx_n_in4),                         //   input,    width = 1,                       .rx_n_in4
		.rx_n_in5                     (hip_serial_rx_n_in5),                         //   input,    width = 1,                       .rx_n_in5
		.rx_n_in6                     (hip_serial_rx_n_in6),                         //   input,    width = 1,                       .rx_n_in6
		.rx_n_in7                     (hip_serial_rx_n_in7),                         //   input,    width = 1,                       .rx_n_in7
		.rx_n_in8                     (hip_serial_rx_n_in8),                         //   input,    width = 1,                       .rx_n_in8
		.rx_n_in9                     (hip_serial_rx_n_in9),                         //   input,    width = 1,                       .rx_n_in9
		.rx_n_in10                    (hip_serial_rx_n_in10),                        //   input,    width = 1,                       .rx_n_in10
		.rx_n_in11                    (hip_serial_rx_n_in11),                        //   input,    width = 1,                       .rx_n_in11
		.rx_n_in12                    (hip_serial_rx_n_in12),                        //   input,    width = 1,                       .rx_n_in12
		.rx_n_in13                    (hip_serial_rx_n_in13),                        //   input,    width = 1,                       .rx_n_in13
		.rx_n_in14                    (hip_serial_rx_n_in14),                        //   input,    width = 1,                       .rx_n_in14
		.rx_n_in15                    (hip_serial_rx_n_in15),                        //   input,    width = 1,                       .rx_n_in15
		.rx_p_in0                     (hip_serial_rx_p_in0),                         //   input,    width = 1,                       .rx_p_in0
		.rx_p_in1                     (hip_serial_rx_p_in1),                         //   input,    width = 1,                       .rx_p_in1
		.rx_p_in2                     (hip_serial_rx_p_in2),                         //   input,    width = 1,                       .rx_p_in2
		.rx_p_in3                     (hip_serial_rx_p_in3),                         //   input,    width = 1,                       .rx_p_in3
		.rx_p_in4                     (hip_serial_rx_p_in4),                         //   input,    width = 1,                       .rx_p_in4
		.rx_p_in5                     (hip_serial_rx_p_in5),                         //   input,    width = 1,                       .rx_p_in5
		.rx_p_in6                     (hip_serial_rx_p_in6),                         //   input,    width = 1,                       .rx_p_in6
		.rx_p_in7                     (hip_serial_rx_p_in7),                         //   input,    width = 1,                       .rx_p_in7
		.rx_p_in8                     (hip_serial_rx_p_in8),                         //   input,    width = 1,                       .rx_p_in8
		.rx_p_in9                     (hip_serial_rx_p_in9),                         //   input,    width = 1,                       .rx_p_in9
		.rx_p_in10                    (hip_serial_rx_p_in10),                        //   input,    width = 1,                       .rx_p_in10
		.rx_p_in11                    (hip_serial_rx_p_in11),                        //   input,    width = 1,                       .rx_p_in11
		.rx_p_in12                    (hip_serial_rx_p_in12),                        //   input,    width = 1,                       .rx_p_in12
		.rx_p_in13                    (hip_serial_rx_p_in13),                        //   input,    width = 1,                       .rx_p_in13
		.rx_p_in14                    (hip_serial_rx_p_in14),                        //   input,    width = 1,                       .rx_p_in14
		.rx_p_in15                    (hip_serial_rx_p_in15),                        //   input,    width = 1,                       .rx_p_in15
		.tx_n_out0                    (hip_serial_tx_n_out0),                        //  output,    width = 1,                       .tx_n_out0
		.tx_n_out1                    (hip_serial_tx_n_out1),                        //  output,    width = 1,                       .tx_n_out1
		.tx_n_out2                    (hip_serial_tx_n_out2),                        //  output,    width = 1,                       .tx_n_out2
		.tx_n_out3                    (hip_serial_tx_n_out3),                        //  output,    width = 1,                       .tx_n_out3
		.tx_n_out4                    (hip_serial_tx_n_out4),                        //  output,    width = 1,                       .tx_n_out4
		.tx_n_out5                    (hip_serial_tx_n_out5),                        //  output,    width = 1,                       .tx_n_out5
		.tx_n_out6                    (hip_serial_tx_n_out6),                        //  output,    width = 1,                       .tx_n_out6
		.tx_n_out7                    (hip_serial_tx_n_out7),                        //  output,    width = 1,                       .tx_n_out7
		.tx_n_out8                    (hip_serial_tx_n_out8),                        //  output,    width = 1,                       .tx_n_out8
		.tx_n_out9                    (hip_serial_tx_n_out9),                        //  output,    width = 1,                       .tx_n_out9
		.tx_n_out10                   (hip_serial_tx_n_out10),                       //  output,    width = 1,                       .tx_n_out10
		.tx_n_out11                   (hip_serial_tx_n_out11),                       //  output,    width = 1,                       .tx_n_out11
		.tx_n_out12                   (hip_serial_tx_n_out12),                       //  output,    width = 1,                       .tx_n_out12
		.tx_n_out13                   (hip_serial_tx_n_out13),                       //  output,    width = 1,                       .tx_n_out13
		.tx_n_out14                   (hip_serial_tx_n_out14),                       //  output,    width = 1,                       .tx_n_out14
		.tx_n_out15                   (hip_serial_tx_n_out15),                       //  output,    width = 1,                       .tx_n_out15
		.tx_p_out0                    (hip_serial_tx_p_out0),                        //  output,    width = 1,                       .tx_p_out0
		.tx_p_out1                    (hip_serial_tx_p_out1),                        //  output,    width = 1,                       .tx_p_out1
		.tx_p_out2                    (hip_serial_tx_p_out2),                        //  output,    width = 1,                       .tx_p_out2
		.tx_p_out3                    (hip_serial_tx_p_out3),                        //  output,    width = 1,                       .tx_p_out3
		.tx_p_out4                    (hip_serial_tx_p_out4),                        //  output,    width = 1,                       .tx_p_out4
		.tx_p_out5                    (hip_serial_tx_p_out5),                        //  output,    width = 1,                       .tx_p_out5
		.tx_p_out6                    (hip_serial_tx_p_out6),                        //  output,    width = 1,                       .tx_p_out6
		.tx_p_out7                    (hip_serial_tx_p_out7),                        //  output,    width = 1,                       .tx_p_out7
		.tx_p_out8                    (hip_serial_tx_p_out8),                        //  output,    width = 1,                       .tx_p_out8
		.tx_p_out9                    (hip_serial_tx_p_out9),                        //  output,    width = 1,                       .tx_p_out9
		.tx_p_out10                   (hip_serial_tx_p_out10),                       //  output,    width = 1,                       .tx_p_out10
		.tx_p_out11                   (hip_serial_tx_p_out11),                       //  output,    width = 1,                       .tx_p_out11
		.tx_p_out12                   (hip_serial_tx_p_out12),                       //  output,    width = 1,                       .tx_p_out12
		.tx_p_out13                   (hip_serial_tx_p_out13),                       //  output,    width = 1,                       .tx_p_out13
		.tx_p_out14                   (hip_serial_tx_p_out14),                       //  output,    width = 1,                       .tx_p_out14
		.tx_p_out15                   (hip_serial_tx_p_out15),                       //  output,    width = 1,                       .tx_p_out15
		.refclk0                      (refclk0_clk),                                 //   input,    width = 1,                refclk0.clk
		.refclk1                      (refclk1_clk),                                 //   input,    width = 1,                refclk1.clk
		.coreclkout_hip               (dut_coreclkout_hip_clk),                      //  output,    width = 1,         coreclkout_hip.clk
		.ninit_done                   (resetip_ninit_done_reset),                    //   input,    width = 1,             ninit_done.reset
		.slow_clk                     (),                                            //  output,    width = 1,               slow_clk.clk
		.pin_perst_n                  (pin_perst_reset_n),                           //   input,    width = 1,              pin_perst.reset_n
		.pin_perst_n_o                ()                                             //  output,    width = 1,          pin_perst_n_o.reset_n
	);
	*/

	pcie_ed_pio0 pio0 (
		.Clk_i                    (dut_coreclkout_hip_clk),                      //   input,     width = 1,              clk.clk
		.Rstn_i                   (dut_p0_reset_status_n_reset),                 //   input,     width = 1,            reset.reset_n
		.pio_clk                  (pio0_pio_master_clk_clk),                     //  output,     width = 1,   pio_master_clk.clk
		.pio_rst_n                (pio0_pio_master_reset_reset),                 //  output,     width = 1, pio_master_reset.reset_n
		.pio_address_o            (pio0_pio_master_address),                     //  output,    width = 64,       pio_master.address
		.pio_read_o               (pio0_pio_master_read),                        //  output,     width = 1,                 .read
		.pio_readdata_i           (pio0_pio_master_readdata),                    //   input,  width = 1024,                 .readdata
		.pio_readdatavalid_i      (pio0_pio_master_readdatavalid),               //   input,     width = 1,                 .readdatavalid
		.pio_write_o              (pio0_pio_master_write),                       //  output,     width = 1,                 .write
		.pio_writedata_o          (pio0_pio_master_writedata),                   //  output,  width = 1024,                 .writedata
		.pio_waitrequest_i        (pio0_pio_master_waitrequest),                 //   input,     width = 1,                 .waitrequest
		.pio_byteenable_o         (pio0_pio_master_byteenable),                  //  output,   width = 128,                 .byteenable
		.pio_response_i           (pio0_pio_master_response),                    //   input,     width = 2,                 .response
		.pio_burstcount_o         (pio0_pio_master_burstcount),                  //  output,     width = 4,                 .burstcount
		.pio_rx_st0_payload_i     (dut_p0_rx_st0_data),                          //   input,   width = 256,       rx_st0_pio.data
		.pio_rx_st0_sop_i         (dut_p0_rx_st0_startofpacket),                 //   input,     width = 1,                 .startofpacket
		.pio_rx_st0_eop_i         (dut_p0_rx_st0_endofpacket),                   //   input,     width = 1,                 .endofpacket
		.pio_rx_st0_dvalid_i      (dut_p0_rx_st0_valid),                         //   input,     width = 1,                 .valid
		.pio_rx_st0_empty_i       (dut_p0_rx_st0_empty),                         //   input,     width = 3,                 .empty
		.pio_rx_st_ready_o        (dut_p0_rx_st0_ready),                         //  output,     width = 1,                 .ready
		.pio_rx_st1_payload_i     (dut_p0_rx_st1_data),                          //   input,   width = 256,       rx_st1_pio.data
		.pio_rx_st1_sop_i         (dut_p0_rx_st1_startofpacket),                 //   input,     width = 1,                 .startofpacket
		.pio_rx_st1_eop_i         (dut_p0_rx_st1_endofpacket),                   //   input,     width = 1,                 .endofpacket
		.pio_rx_st1_dvalid_i      (dut_p0_rx_st1_valid),                         //   input,     width = 1,                 .valid
		.pio_rx_st1_empty_i       (dut_p0_rx_st1_empty),                         //   input,     width = 3,                 .empty
		.pio_rx_st2_payload_i     (dut_p0_rx_st2_data),                          //   input,   width = 256,       rx_st2_pio.data
		.pio_rx_st2_sop_i         (dut_p0_rx_st2_startofpacket),                 //   input,     width = 1,                 .startofpacket
		.pio_rx_st2_eop_i         (dut_p0_rx_st2_endofpacket),                   //   input,     width = 1,                 .endofpacket
		.pio_rx_st2_dvalid_i      (dut_p0_rx_st2_valid),                         //   input,     width = 1,                 .valid
		.pio_rx_st2_empty_i       (dut_p0_rx_st2_empty),                         //   input,     width = 3,                 .empty
		.pio_rx_st3_payload_i     (dut_p0_rx_st3_data),                          //   input,   width = 256,       rx_st3_pio.data
		.pio_rx_st3_sop_i         (dut_p0_rx_st3_startofpacket),                 //   input,     width = 1,                 .startofpacket
		.pio_rx_st3_eop_i         (dut_p0_rx_st3_endofpacket),                   //   input,     width = 1,                 .endofpacket
		.pio_rx_st3_dvalid_i      (dut_p0_rx_st3_valid),                         //   input,     width = 1,                 .valid
		.pio_rx_st3_empty_i       (dut_p0_rx_st3_empty),                         //   input,     width = 3,                 .empty
		.rx_st_hcrdt_init_o       (pio0_rx_st0_pio_misc_rx_st_hcrdt_init),       //  output,     width = 3,  rx_st0_pio_misc.rx_st_Hcrdt_init
		.rx_st_hcrdt_update_o     (pio0_rx_st0_pio_misc_rx_st_hcrdt_update),     //  output,     width = 3,                 .rx_st_Hcrdt_update
		.rx_st_hcrdt_update_cnt_o (pio0_rx_st0_pio_misc_rx_st_hcrdt_update_cnt), //  output,     width = 6,                 .rx_st_Hcrdt_update_cnt
		.rx_st_hcrdt_init_ack_i   (dut_p0_rx_st_misc_rx_st_hcrdt_init_ack),      //   input,     width = 3,                 .rx_st_Hcrdt_init_ack
		.rx_st_dcrdt_init_o       (pio0_rx_st0_pio_misc_rx_st_dcrdt_init),       //  output,     width = 3,                 .rx_st_Dcrdt_init
		.rx_st_dcrdt_update_o     (pio0_rx_st0_pio_misc_rx_st_dcrdt_update),     //  output,     width = 3,                 .rx_st_Dcrdt_update
		.rx_st_dcrdt_update_cnt_o (pio0_rx_st0_pio_misc_rx_st_dcrdt_update_cnt), //  output,    width = 12,                 .rx_st_Dcrdt_update_cnt
		.rx_st_dcrdt_init_ack_i   (dut_p0_rx_st_misc_rx_st_dcrdt_init_ack),      //   input,     width = 3,                 .rx_st_Dcrdt_init_ack
		.pio_rx_st0_header_i      (dut_p0_rx_st_misc_rx_st0_hdr),                //   input,   width = 128,                 .rx_st0_hdr
		.pio_rx_st0_tlp_prfx_i    (dut_p0_rx_st_misc_rx_st0_prefix),             //   input,    width = 32,                 .rx_st0_prefix
		.pio_rx_st0_hvalid_i      (dut_p0_rx_st_misc_rx_st0_hvalid),             //   input,     width = 1,                 .rx_st0_hvalid
		.pio_rx_st0_pvalid_i      (dut_p0_rx_st_misc_rx_st0_pvalid),             //   input,     width = 1,                 .rx_st0_pvalid
		.pio_rx_st0_bar_i         (dut_p0_rx_st_misc_rx_st0_bar),                //   input,     width = 3,                 .rx_st0_bar
		.pio_rx_st1_header_i      (dut_p0_rx_st_misc_rx_st1_hdr),                //   input,   width = 128,                 .rx_st1_hdr
		.pio_rx_st1_tlp_prfx_i    (dut_p0_rx_st_misc_rx_st1_prefix),             //   input,    width = 32,                 .rx_st1_prefix
		.pio_rx_st1_hvalid_i      (dut_p0_rx_st_misc_rx_st1_hvalid),             //   input,     width = 1,                 .rx_st1_hvalid
		.pio_rx_st1_pvalid_i      (dut_p0_rx_st_misc_rx_st1_pvalid),             //   input,     width = 1,                 .rx_st1_pvalid
		.pio_rx_st1_bar_i         (dut_p0_rx_st_misc_rx_st1_bar),                //   input,     width = 3,                 .rx_st1_bar
		.pio_rx_st2_header_i      (dut_p0_rx_st_misc_rx_st2_hdr),                //   input,   width = 128,                 .rx_st2_hdr
		.pio_rx_st2_tlp_prfx_i    (dut_p0_rx_st_misc_rx_st2_prefix),             //   input,    width = 32,                 .rx_st2_prefix
		.pio_rx_st2_hvalid_i      (dut_p0_rx_st_misc_rx_st2_hvalid),             //   input,     width = 1,                 .rx_st2_hvalid
		.pio_rx_st2_pvalid_i      (dut_p0_rx_st_misc_rx_st2_pvalid),             //   input,     width = 1,                 .rx_st2_pvalid
		.pio_rx_st2_bar_i         (dut_p0_rx_st_misc_rx_st2_bar),                //   input,     width = 3,                 .rx_st2_bar
		.pio_rx_st3_header_i      (dut_p0_rx_st_misc_rx_st3_hdr),                //   input,   width = 128,                 .rx_st3_hdr
		.pio_rx_st3_tlp_prfx_i    (dut_p0_rx_st_misc_rx_st3_prefix),             //   input,    width = 32,                 .rx_st3_prefix
		.pio_rx_st3_hvalid_i      (dut_p0_rx_st_misc_rx_st3_hvalid),             //   input,     width = 1,                 .rx_st3_hvalid
		.pio_rx_st3_pvalid_i      (dut_p0_rx_st_misc_rx_st3_pvalid),             //   input,     width = 1,                 .rx_st3_pvalid
		.pio_rx_st3_bar_i         (dut_p0_rx_st_misc_rx_st3_bar),                //   input,     width = 3,                 .rx_st3_bar
		.pio_tx_st0_payload_o     (pio0_tx_st0_pio_data),                        //  output,   width = 256,       tx_st0_pio.data
		.pio_tx_st0_sop_o         (pio0_tx_st0_pio_startofpacket),               //  output,     width = 1,                 .startofpacket
		.pio_tx_st0_eop_o         (pio0_tx_st0_pio_endofpacket),                 //  output,     width = 1,                 .endofpacket
		.pio_tx_st0_dvalid_o      (pio0_tx_st0_pio_valid),                       //  output,     width = 1,                 .valid
		.pio_tx_st_ready_i        (pio0_tx_st0_pio_ready),                       //   input,     width = 1,                 .ready
		.pio_tx_st1_payload_o     (pio0_tx_st1_pio_data),                        //  output,   width = 256,       tx_st1_pio.data
		.pio_tx_st1_sop_o         (pio0_tx_st1_pio_startofpacket),               //  output,     width = 1,                 .startofpacket
		.pio_tx_st1_eop_o         (pio0_tx_st1_pio_endofpacket),                 //  output,     width = 1,                 .endofpacket
		.pio_tx_st1_dvalid_o      (pio0_tx_st1_pio_valid),                       //  output,     width = 1,                 .valid
		.pio_tx_st2_payload_o     (pio0_tx_st2_pio_data),                        //  output,   width = 256,       tx_st2_pio.data
		.pio_tx_st2_sop_o         (pio0_tx_st2_pio_startofpacket),               //  output,     width = 1,                 .startofpacket
		.pio_tx_st2_eop_o         (pio0_tx_st2_pio_endofpacket),                 //  output,     width = 1,                 .endofpacket
		.pio_tx_st2_dvalid_o      (pio0_tx_st2_pio_valid),                       //  output,     width = 1,                 .valid
		.pio_tx_st3_payload_o     (pio0_tx_st3_pio_data),                        //  output,   width = 256,       tx_st3_pio.data
		.pio_tx_st3_sop_o         (pio0_tx_st3_pio_startofpacket),               //  output,     width = 1,                 .startofpacket
		.pio_tx_st3_eop_o         (pio0_tx_st3_pio_endofpacket),                 //  output,     width = 1,                 .endofpacket
		.pio_tx_st3_dvalid_o      (pio0_tx_st3_pio_valid),                       //  output,     width = 1,                 .valid
		.pio_tx_st0_header_o      (pio0_tx_st0_pio_misc_tx_st0_hdr),             //  output,   width = 128,  tx_st0_pio_misc.tx_st0_hdr
		.pio_tx_st1_header_o      (pio0_tx_st0_pio_misc_tx_st1_hdr),             //  output,   width = 128,                 .tx_st1_hdr
		.pio_tx_st2_header_o      (pio0_tx_st0_pio_misc_tx_st2_hdr),             //  output,   width = 128,                 .tx_st2_hdr
		.pio_tx_st3_header_o      (pio0_tx_st0_pio_misc_tx_st3_hdr),             //  output,   width = 128,                 .tx_st3_hdr
		.tx_st_hcrdt_init_i       (dut_p0_tx_st_misc_tx_st_hcrdt_init),          //   input,     width = 3,                 .tx_st_Hcrdt_init
		.tx_st_hcrdt_update_i     (dut_p0_tx_st_misc_tx_st_hcrdt_update),        //   input,     width = 3,                 .tx_st_Hcrdt_update
		.tx_st_hcrdt_update_cnt_i (dut_p0_tx_st_misc_tx_st_hcrdt_update_cnt),    //   input,     width = 6,                 .tx_st_Hcrdt_update_cnt
		.tx_st_hcrdt_init_ack_o   (pio0_tx_st0_pio_misc_tx_st_hcrdtt_init_ack),  //  output,     width = 3,                 .tx_st_Hcrdtt_init_ack
		.tx_st_dcrdt_init_i       (dut_p0_tx_st_misc_tx_st_dcrdt_init),          //   input,     width = 3,                 .tx_st_Dcrdt_init
		.tx_st_dcrdt_update_i     (dut_p0_tx_st_misc_tx_st_dcrdt_update),        //   input,     width = 3,                 .tx_st_Dcrdt_update
		.tx_st_dcrdt_update_cnt_i (dut_p0_tx_st_misc_tx_st_dcrdt_update_cnt),    //   input,    width = 12,                 .tx_st_Dcrdt_update_cnt
		.tx_st_dcrdt_init_ack_o   (pio0_tx_st0_pio_misc_tx_st_dcrdt_init_ack),   //  output,     width = 3,                 .tx_st_Dcrdt_init_ack
		.pio_tx_st0_prefix_o      (pio0_tx_st0_pio_misc_tx_st0_prefix),          //  output,    width = 32,                 .tx_st0_prefix
		.pio_tx_st0_hvalid_o      (pio0_tx_st0_pio_misc_tx_st0_hvalid),          //  output,     width = 1,                 .tx_st0_hvalid
		.pio_tx_st0_pvalid_o      (pio0_tx_st0_pio_misc_tx_st0_pvalid),          //  output,     width = 1,                 .tx_st0_pvalid
		.pio_tx_st1_prefix_o      (pio0_tx_st0_pio_misc_tx_st1_prefix),          //  output,    width = 32,                 .tx_st1_prefix
		.pio_tx_st1_hvalid_o      (pio0_tx_st0_pio_misc_tx_st1_hvalid),          //  output,     width = 1,                 .tx_st1_hvalid
		.pio_tx_st1_pvalid_o      (pio0_tx_st0_pio_misc_tx_st1_pvalid),          //  output,     width = 1,                 .tx_st1_pvalid
		.pio_tx_st2_prefix_o      (pio0_tx_st0_pio_misc_tx_st2_prefix),          //  output,    width = 32,                 .tx_st2_prefix
		.pio_tx_st2_hvalid_o      (pio0_tx_st0_pio_misc_tx_st2_hvalid),          //  output,     width = 1,                 .tx_st2_hvalid
		.pio_tx_st2_pvalid_o      (pio0_tx_st0_pio_misc_tx_st2_pvalid),          //  output,     width = 1,                 .tx_st2_pvalid
		.pio_tx_st3_prefix_o      (pio0_tx_st0_pio_misc_tx_st3_prefix),          //  output,    width = 32,                 .tx_st3_prefix
		.pio_tx_st3_hvalid_o      (pio0_tx_st0_pio_misc_tx_st3_hvalid),          //  output,     width = 1,                 .tx_st3_hvalid
		.pio_tx_st3_pvalid_o      (pio0_tx_st0_pio_misc_tx_st3_pvalid)           //  output,     width = 1,                 .tx_st3_pvalid
	);

	/*
	pcie_ed_resetIP resetip (
		.ninit_done (resetip_ninit_done_reset)  //  output,  width = 1, ninit_done.reset
	);
	*/

	pcie_ed_altera_mm_interconnect_1920_sx2feoa mm_interconnect_0 (
		.pio0_pio_master_address                                      (pio0_pio_master_address),              //   input,    width = 64,                                        pio0_pio_master.address
		.pio0_pio_master_waitrequest                                  (pio0_pio_master_waitrequest),          //  output,     width = 1,                                                       .waitrequest
		.pio0_pio_master_burstcount                                   (pio0_pio_master_burstcount),           //   input,     width = 4,                                                       .burstcount
		.pio0_pio_master_byteenable                                   (pio0_pio_master_byteenable),           //   input,   width = 128,                                                       .byteenable
		.pio0_pio_master_read                                         (pio0_pio_master_read),                 //   input,     width = 1,                                                       .read
		.pio0_pio_master_readdata                                     (pio0_pio_master_readdata),             //  output,  width = 1024,                                                       .readdata
		.pio0_pio_master_readdatavalid                                (pio0_pio_master_readdatavalid),        //  output,     width = 1,                                                       .readdatavalid
		.pio0_pio_master_write                                        (pio0_pio_master_write),                //   input,     width = 1,                                                       .write
		.pio0_pio_master_writedata                                    (pio0_pio_master_writedata),            //   input,  width = 1024,                                                       .writedata
		.pio0_pio_master_response                                     (pio0_pio_master_response),             //  output,     width = 2,                                                       .response
		.MEM0_s1_address                                              (mm_interconnect_0_mem0_s1_address),    //  output,     width = 8,                                                MEM0_s1.address
		.MEM0_s1_write                                                (mm_interconnect_0_mem0_s1_write),      //  output,     width = 1,                                                       .write
		.MEM0_s1_readdata                                             (mm_interconnect_0_mem0_s1_readdata),   //   input,  width = 1024,                                                       .readdata
		.MEM0_s1_writedata                                            (mm_interconnect_0_mem0_s1_writedata),  //  output,  width = 1024,                                                       .writedata
		.MEM0_s1_byteenable                                           (mm_interconnect_0_mem0_s1_byteenable), //  output,   width = 128,                                                       .byteenable
		.MEM0_s1_chipselect                                           (mm_interconnect_0_mem0_s1_chipselect), //  output,     width = 1,                                                       .chipselect
		.MEM0_s1_clken                                                (mm_interconnect_0_mem0_s1_clken),      //  output,     width = 1,                                                       .clken
		.MEM0_reset1_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),       //   input,     width = 1,                      MEM0_reset1_reset_bridge_in_reset.reset
		.pio0_pio_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),       //   input,     width = 1, pio0_pio_master_translator_reset_reset_bridge_in_reset.reset
		.pio0_pio_master_clk_clk                                      (pio0_pio_master_clk_clk)               //   input,     width = 1,                                    pio0_pio_master_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pio0_pio_master_reset_reset),   //   input,  width = 1, reset_in0.reset
		.clk            (pio0_pio_master_clk_clk),        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "5SOp2wqjkMCvRs5H/8cuggoPFnOYOVi/4/bu0Ttyg6RGDyAtuEiXM6zkpXTknpEbjlGv1qJhvF6QsriNG9ARPZ7JmiU3BFWTE9LqHzcFT7tPdS7N8boITkYqxt5v97iIEFF1Inp38Z2ZjsNVDWx8i62p0LDZ9g0btA81KMjFRSEqWO+7zoj3fGDFVT4C92nEu4HzJ3Vn/6UckyxLHS+UBqQ5vFQM1/jRM3utVd+aJiI9FU0P85IKaz4+z6nlGkM6QzRwJ1WwrGsqWNSMNQvF85qa6woc5NJpAyP+OIY0K4YoS04zrKEiFe/1AAWhfgbHi6CrYCJscUwuJ1QpSYtxXwce1zBRr0GDmzQCGYOHhhZrifeG6gxoDJvst1a8ix8XFxGFVY3qSs7gHoxHX394JBx2WatL4sVxPRuQFkA7Ekw5fc8LXKqEHcGw0C15jdQfudUn4whkIIaW0wSYBVgBkGey/5MkjDFd6A+oFvVVKK93lG/e389/R1qdwFV0BhPIML2E0prd65vf3np0Vy1XJvooJ9pw0/bGTNq03QlpE+XBluRnQdK4MS89zs3rkxMN/Tu2eviOaLHKw7KFIvlwKXGip878ly8wirpVFPW+uxoUS2RJmaVpu6tPvovzKsTdqsW+RyTi8fqHjyAZUzo2/vOpFQEFul9sNHgzBIyCOfIu9Ek0UHIcNUMO7zSxXq5xV0MnOGiHJJLIwuiRlRUAbrKintHecROeXPI/8ty/QXIN0z+oz07H8cJ0NV+tdHnT1cJTXvgtlINNF/qf2uc8jovgkM4/poijuoYiZ9ZOPbDAv3h2OE+elp1X3YNCa3JLLo8azIvJe4KxwVrAv6Vn4ptCcpQ3Uy+q1tmUb4WjRO1zwUmeX6i2J09uBZ6j4qLYrr6IqDSsO6VuhRC2hxwByN97mPYpPN/5GbtYyqqy3jAd99QES8j+bED87kmmQVSWKPQ8BPu3sBnmXv4J41l6ZY1lTzSwdHTDKLnX9IIZkpXDiXGqsIVrbZtaEYJeq08n"
`endif